library verilog;
use verilog.vl_types.all;
entity tb_top_npu_system is
end tb_top_npu_system;
