library verilog;
use verilog.vl_types.all;
entity EMCU is
    port(
        FCLK            : in     vl_logic;
        PORESETN        : in     vl_logic;
        SYSRESETN       : in     vl_logic;
        RTCSRCCLK       : in     vl_logic;
        IOEXPOUTPUTO    : out    vl_logic_vector(15 downto 0);
        IOEXPOUTPUTENO  : out    vl_logic_vector(15 downto 0);
        IOEXPINPUTI     : in     vl_logic_vector(15 downto 0);
        UART0TXDO       : out    vl_logic;
        UART1TXDO       : out    vl_logic;
        UART0BAUDTICK   : out    vl_logic;
        UART1BAUDTICK   : out    vl_logic;
        UART0RXDI       : in     vl_logic;
        UART1RXDI       : in     vl_logic;
        INTMONITOR      : out    vl_logic;
        MTXHRESETN      : out    vl_logic;
        SRAM0ADDR       : out    vl_logic_vector(12 downto 0);
        SRAM0WREN       : out    vl_logic_vector(3 downto 0);
        SRAM0WDATA      : out    vl_logic_vector(31 downto 0);
        SRAM0CS         : out    vl_logic;
        SRAM0RDATA      : in     vl_logic_vector(31 downto 0);
        TARGFLASH0HSEL  : out    vl_logic;
        TARGFLASH0HADDR : out    vl_logic_vector(28 downto 0);
        TARGFLASH0HTRANS: out    vl_logic_vector(1 downto 0);
        TARGFLASH0HSIZE : out    vl_logic_vector(2 downto 0);
        TARGFLASH0HBURST: out    vl_logic_vector(2 downto 0);
        TARGFLASH0HREADYMUX: out    vl_logic;
        TARGFLASH0HRDATA: in     vl_logic_vector(31 downto 0);
        TARGFLASH0HRUSER: in     vl_logic_vector(2 downto 0);
        TARGFLASH0HRESP : in     vl_logic;
        TARGFLASH0EXRESP: in     vl_logic;
        TARGFLASH0HREADYOUT: in     vl_logic;
        TARGEXP0HSEL    : out    vl_logic;
        TARGEXP0HADDR   : out    vl_logic_vector(31 downto 0);
        TARGEXP0HTRANS  : out    vl_logic_vector(1 downto 0);
        TARGEXP0HWRITE  : out    vl_logic;
        TARGEXP0HSIZE   : out    vl_logic_vector(2 downto 0);
        TARGEXP0HBURST  : out    vl_logic_vector(2 downto 0);
        TARGEXP0HPROT   : out    vl_logic_vector(3 downto 0);
        TARGEXP0MEMATTR : out    vl_logic_vector(1 downto 0);
        TARGEXP0EXREQ   : out    vl_logic;
        TARGEXP0HMASTER : out    vl_logic_vector(3 downto 0);
        TARGEXP0HWDATA  : out    vl_logic_vector(31 downto 0);
        TARGEXP0HMASTLOCK: out    vl_logic;
        TARGEXP0HREADYMUX: out    vl_logic;
        TARGEXP0HAUSER  : out    vl_logic;
        TARGEXP0HWUSER  : out    vl_logic_vector(3 downto 0);
        TARGEXP0HRDATA  : in     vl_logic_vector(31 downto 0);
        TARGEXP0HREADYOUT: in     vl_logic;
        TARGEXP0HRESP   : in     vl_logic;
        TARGEXP0EXRESP  : in     vl_logic;
        TARGEXP0HRUSER  : in     vl_logic_vector(2 downto 0);
        INITEXP0HRDATA  : out    vl_logic_vector(31 downto 0);
        INITEXP0HREADY  : out    vl_logic;
        INITEXP0HRESP   : out    vl_logic;
        INITEXP0EXRESP  : out    vl_logic;
        INITEXP0HRUSER  : out    vl_logic_vector(2 downto 0);
        INITEXP0HSEL    : in     vl_logic;
        INITEXP0HADDR   : in     vl_logic_vector(31 downto 0);
        INITEXP0HTRANS  : in     vl_logic_vector(1 downto 0);
        INITEXP0HWRITE  : in     vl_logic;
        INITEXP0HSIZE   : in     vl_logic_vector(2 downto 0);
        INITEXP0HBURST  : in     vl_logic_vector(2 downto 0);
        INITEXP0HPROT   : in     vl_logic_vector(3 downto 0);
        INITEXP0MEMATTR : in     vl_logic_vector(1 downto 0);
        INITEXP0EXREQ   : in     vl_logic;
        INITEXP0HMASTER : in     vl_logic_vector(3 downto 0);
        INITEXP0HWDATA  : in     vl_logic_vector(31 downto 0);
        INITEXP0HMASTLOCK: in     vl_logic;
        INITEXP0HAUSER  : in     vl_logic;
        INITEXP0HWUSER  : in     vl_logic_vector(3 downto 0);
        APBTARGEXP2PSTRB: out    vl_logic_vector(3 downto 0);
        APBTARGEXP2PPROT: out    vl_logic_vector(2 downto 0);
        APBTARGEXP2PSEL : out    vl_logic;
        APBTARGEXP2PENABLE: out    vl_logic;
        APBTARGEXP2PADDR: out    vl_logic_vector(11 downto 0);
        APBTARGEXP2PWRITE: out    vl_logic;
        APBTARGEXP2PWDATA: out    vl_logic_vector(31 downto 0);
        APBTARGEXP2PRDATA: in     vl_logic_vector(31 downto 0);
        APBTARGEXP2PREADY: in     vl_logic;
        APBTARGEXP2PSLVERR: in     vl_logic;
        MTXREMAP        : in     vl_logic_vector(3 downto 0);
        DAPTDO          : out    vl_logic;
        DAPJTAGNSW      : out    vl_logic;
        DAPNTDOEN       : out    vl_logic;
        DAPSWDITMS      : in     vl_logic;
        DAPTDI          : in     vl_logic;
        DAPNTRST        : in     vl_logic;
        DAPSWCLKTCK     : in     vl_logic;
        TPIUTRACEDATA   : out    vl_logic_vector(3 downto 0);
        TPIUTRACECLK    : out    vl_logic;
        GPINT           : in     vl_logic_vector(4 downto 0);
        FLASHERR        : in     vl_logic;
        FLASHINT        : in     vl_logic
    );
end EMCU;
