library verilog;
use verilog.vl_types.all;
entity BANDGAP is
    port(
        BGEN            : in     vl_logic
    );
end BANDGAP;
