library verilog;
use verilog.vl_types.all;
entity rPLL is
    generic(
        FCLKIN          : string  := "100.0";
        DYN_IDIV_SEL    : string  := "false";
        IDIV_SEL        : integer := 0;
        DYN_FBDIV_SEL   : string  := "false";
        FBDIV_SEL       : integer := 0;
        DYN_ODIV_SEL    : string  := "false";
        ODIV_SEL        : integer := 8;
        PSDA_SEL        : string  := "0000";
        DYN_DA_EN       : string  := "false";
        DUTYDA_SEL      : string  := "1000";
        CLKOUT_FT_DIR   : vl_logic := Hi1;
        CLKOUTP_FT_DIR  : vl_logic := Hi1;
        CLKOUT_DLY_STEP : integer := 0;
        CLKOUTP_DLY_STEP: integer := 0;
        CLKFB_SEL       : string  := "internal";
        CLKOUT_BYPASS   : string  := "false";
        CLKOUTP_BYPASS  : string  := "false";
        CLKOUTD_BYPASS  : string  := "false";
        DYN_SDIV_SEL    : integer := 2;
        CLKOUTD_SRC     : string  := "CLKOUT";
        CLKOUTD3_SRC    : string  := "CLKOUT";
        DEVICE          : string  := "GW1N-4"
    );
    port(
        CLKOUT          : out    vl_logic;
        CLKOUTP         : out    vl_logic;
        CLKOUTD         : out    vl_logic;
        CLKOUTD3        : out    vl_logic;
        LOCK            : out    vl_logic;
        CLKIN           : in     vl_logic;
        CLKFB           : in     vl_logic;
        FBDSEL          : in     vl_logic_vector(5 downto 0);
        IDSEL           : in     vl_logic_vector(5 downto 0);
        ODSEL           : in     vl_logic_vector(5 downto 0);
        DUTYDA          : in     vl_logic_vector(3 downto 0);
        PSDA            : in     vl_logic_vector(3 downto 0);
        FDLY            : in     vl_logic_vector(3 downto 0);
        RESET           : in     vl_logic;
        RESET_P         : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of FCLKIN : constant is 1;
    attribute mti_svvh_generic_type of DYN_IDIV_SEL : constant is 1;
    attribute mti_svvh_generic_type of IDIV_SEL : constant is 1;
    attribute mti_svvh_generic_type of DYN_FBDIV_SEL : constant is 1;
    attribute mti_svvh_generic_type of FBDIV_SEL : constant is 1;
    attribute mti_svvh_generic_type of DYN_ODIV_SEL : constant is 1;
    attribute mti_svvh_generic_type of ODIV_SEL : constant is 1;
    attribute mti_svvh_generic_type of PSDA_SEL : constant is 1;
    attribute mti_svvh_generic_type of DYN_DA_EN : constant is 1;
    attribute mti_svvh_generic_type of DUTYDA_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT_FT_DIR : constant is 1;
    attribute mti_svvh_generic_type of CLKOUTP_FT_DIR : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT_DLY_STEP : constant is 1;
    attribute mti_svvh_generic_type of CLKOUTP_DLY_STEP : constant is 1;
    attribute mti_svvh_generic_type of CLKFB_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT_BYPASS : constant is 1;
    attribute mti_svvh_generic_type of CLKOUTP_BYPASS : constant is 1;
    attribute mti_svvh_generic_type of CLKOUTD_BYPASS : constant is 1;
    attribute mti_svvh_generic_type of DYN_SDIV_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKOUTD_SRC : constant is 1;
    attribute mti_svvh_generic_type of CLKOUTD3_SRC : constant is 1;
    attribute mti_svvh_generic_type of DEVICE : constant is 1;
end rPLL;
