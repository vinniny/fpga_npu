library verilog;
use verilog.vl_types.all;
entity tb_spi_slave is
end tb_spi_slave;
