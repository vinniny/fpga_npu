library verilog;
use verilog.vl_types.all;
entity PWRGRD is
    port(
        PDEN            : in     vl_logic
    );
end PWRGRD;
