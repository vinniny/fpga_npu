library verilog;
use verilog.vl_types.all;
entity IDES16 is
    generic(
        GSREN           : string  := "false";
        LSREN           : string  := "true"
    );
    port(
        Q0              : out    vl_logic;
        Q1              : out    vl_logic;
        Q2              : out    vl_logic;
        Q3              : out    vl_logic;
        Q4              : out    vl_logic;
        Q5              : out    vl_logic;
        Q6              : out    vl_logic;
        Q7              : out    vl_logic;
        Q8              : out    vl_logic;
        Q9              : out    vl_logic;
        Q10             : out    vl_logic;
        Q11             : out    vl_logic;
        Q12             : out    vl_logic;
        Q13             : out    vl_logic;
        Q14             : out    vl_logic;
        Q15             : out    vl_logic;
        D               : in     vl_logic;
        CALIB           : in     vl_logic;
        PCLK            : in     vl_logic;
        FCLK            : in     vl_logic;
        RESET           : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of GSREN : constant is 1;
    attribute mti_svvh_generic_type of LSREN : constant is 1;
end IDES16;
