library verilog;
use verilog.vl_types.all;
entity tb_gowin_multaddalu is
end tb_gowin_multaddalu;
