library verilog;
use verilog.vl_types.all;
entity tb_sram_A is
end tb_sram_A;
