library verilog;
use verilog.vl_types.all;
entity tb_matrix_convolution_debug is
end tb_matrix_convolution_debug;
