library verilog;
use verilog.vl_types.all;
entity tb_sram_B is
end tb_sram_B;
