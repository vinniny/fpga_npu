library verilog;
use verilog.vl_types.all;
entity tb_sram_C is
end tb_sram_C;
