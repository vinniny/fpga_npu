library verilog;
use verilog.vl_types.all;
entity VCC is
    port(
        V               : out    vl_logic
    );
end VCC;
