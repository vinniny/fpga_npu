library verilog;
use verilog.vl_types.all;
entity tb_tile_processor is
end tb_tile_processor;
