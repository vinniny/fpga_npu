library verilog;
use verilog.vl_types.all;
entity MIPI_DPHY_RX is
    generic(
        ALIGN_BYTE      : vl_logic_vector(0 to 7) := (Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0);
        MIPI_LANE0_EN   : vl_logic := Hi0;
        MIPI_LANE1_EN   : vl_logic := Hi0;
        MIPI_LANE2_EN   : vl_logic := Hi0;
        MIPI_LANE3_EN   : vl_logic := Hi0;
        MIPI_CK_EN      : vl_logic := Hi1;
        SYNC_CLK_SEL    : vl_logic := Hi0
    );
    port(
        D0LN_HSRXD      : out    vl_logic_vector(15 downto 0);
        D1LN_HSRXD      : out    vl_logic_vector(15 downto 0);
        D2LN_HSRXD      : out    vl_logic_vector(15 downto 0);
        D3LN_HSRXD      : out    vl_logic_vector(15 downto 0);
        D0LN_HSRXD_VLD  : out    vl_logic;
        D1LN_HSRXD_VLD  : out    vl_logic;
        D2LN_HSRXD_VLD  : out    vl_logic;
        D3LN_HSRXD_VLD  : out    vl_logic;
        DI_LPRX0_N      : out    vl_logic;
        DI_LPRX0_P      : out    vl_logic;
        DI_LPRX1_N      : out    vl_logic;
        DI_LPRX1_P      : out    vl_logic;
        DI_LPRX2_N      : out    vl_logic;
        DI_LPRX2_P      : out    vl_logic;
        DI_LPRX3_N      : out    vl_logic;
        DI_LPRX3_P      : out    vl_logic;
        DI_LPRXCK_N     : out    vl_logic;
        DI_LPRXCK_P     : out    vl_logic;
        RX_CLK_O        : out    vl_logic;
        DESKEW_ERROR    : out    vl_logic;
        CK_N            : inout  vl_logic;
        CK_P            : inout  vl_logic;
        RX0_N           : inout  vl_logic;
        RX0_P           : inout  vl_logic;
        RX1_N           : inout  vl_logic;
        RX1_P           : inout  vl_logic;
        RX2_N           : inout  vl_logic;
        RX2_P           : inout  vl_logic;
        RX3_N           : inout  vl_logic;
        RX3_P           : inout  vl_logic;
        LPRX_EN_CK      : in     vl_logic;
        LPRX_EN_D0      : in     vl_logic;
        LPRX_EN_D1      : in     vl_logic;
        LPRX_EN_D2      : in     vl_logic;
        LPRX_EN_D3      : in     vl_logic;
        HSRX_ODTEN_CK   : in     vl_logic;
        HSRX_ODTEN_D0   : in     vl_logic;
        HSRX_ODTEN_D1   : in     vl_logic;
        HSRX_ODTEN_D2   : in     vl_logic;
        HSRX_ODTEN_D3   : in     vl_logic;
        D0LN_HSRX_DREN  : in     vl_logic;
        D1LN_HSRX_DREN  : in     vl_logic;
        D2LN_HSRX_DREN  : in     vl_logic;
        D3LN_HSRX_DREN  : in     vl_logic;
        HSRX_EN_CK      : in     vl_logic;
        DESKEW_REQ      : in     vl_logic;
        HS_8BIT_MODE    : in     vl_logic;
        RX_CLK_1X       : in     vl_logic;
        RX_INVERT       : in     vl_logic;
        LALIGN_EN       : in     vl_logic;
        WALIGN_BY       : in     vl_logic;
        DO_LPTX0_N      : in     vl_logic;
        DO_LPTX0_P      : in     vl_logic;
        DO_LPTX1_N      : in     vl_logic;
        DO_LPTX1_P      : in     vl_logic;
        DO_LPTX2_N      : in     vl_logic;
        DO_LPTX2_P      : in     vl_logic;
        DO_LPTX3_N      : in     vl_logic;
        DO_LPTX3_P      : in     vl_logic;
        DO_LPTXCK_N     : in     vl_logic;
        DO_LPTXCK_P     : in     vl_logic;
        LPTX_EN_CK      : in     vl_logic;
        LPTX_EN_D0      : in     vl_logic;
        LPTX_EN_D1      : in     vl_logic;
        LPTX_EN_D2      : in     vl_logic;
        LPTX_EN_D3      : in     vl_logic;
        BYTE_LENDIAN    : in     vl_logic;
        HSRX_STOP       : in     vl_logic;
        LPRX_ULP_LN0    : in     vl_logic;
        LPRX_ULP_LN1    : in     vl_logic;
        LPRX_ULP_LN2    : in     vl_logic;
        LPRX_ULP_LN3    : in     vl_logic;
        LPRX_ULP_CK     : in     vl_logic;
        PWRON           : in     vl_logic;
        RESET           : in     vl_logic;
        DESKEW_LNSEL    : in     vl_logic_vector(2 downto 0);
        DESKEW_MTH      : in     vl_logic_vector(7 downto 0);
        DESKEW_OWVAL    : in     vl_logic_vector(6 downto 0);
        DRST_N          : in     vl_logic;
        ONE_BYTE0_MATCH : in     vl_logic;
        WORD_LENDIAN    : in     vl_logic;
        FIFO_RD_STD     : in     vl_logic_vector(2 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of ALIGN_BYTE : constant is 1;
    attribute mti_svvh_generic_type of MIPI_LANE0_EN : constant is 1;
    attribute mti_svvh_generic_type of MIPI_LANE1_EN : constant is 1;
    attribute mti_svvh_generic_type of MIPI_LANE2_EN : constant is 1;
    attribute mti_svvh_generic_type of MIPI_LANE3_EN : constant is 1;
    attribute mti_svvh_generic_type of MIPI_CK_EN : constant is 1;
    attribute mti_svvh_generic_type of SYNC_CLK_SEL : constant is 1;
end MIPI_DPHY_RX;
