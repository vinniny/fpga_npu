library verilog;
use verilog.vl_types.all;
entity GSR is
    port(
        GSRI            : in     vl_logic
    );
end GSR;
