library verilog;
use verilog.vl_types.all;
entity tb_matrix_dot is
end tb_matrix_dot;
