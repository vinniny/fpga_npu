library verilog;
use verilog.vl_types.all;
entity tb_matrix_multiplier is
end tb_matrix_multiplier;
