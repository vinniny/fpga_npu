library verilog;
use verilog.vl_types.all;
entity tb_gowin_rpll is
end tb_gowin_rpll;
