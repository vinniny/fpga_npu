library verilog;
use verilog.vl_types.all;
entity BUFS is
    port(
        O               : out    vl_logic;
        I               : in     vl_logic
    );
end BUFS;
