library verilog;
use verilog.vl_types.all;
entity PLLO is
    generic(
        FCLKIN          : string  := "100.0";
        DYN_IDIV_SEL    : string  := "FALSE";
        IDIV_SEL        : integer := 0;
        DYN_FBDIV_SEL   : string  := "FALSE";
        FBDIV_SEL       : integer := 0;
        DYN_ODIVA_SEL   : string  := "FALSE";
        ODIVA_SEL       : integer := 6;
        DYN_ODIVB_SEL   : string  := "FALSE";
        ODIVB_SEL       : integer := 6;
        DYN_ODIVC_SEL   : string  := "FALSE";
        ODIVC_SEL       : integer := 6;
        DYN_ODIVD_SEL   : string  := "FALSE";
        ODIVD_SEL       : integer := 6;
        CLKOUTA_EN      : string  := "TRUE";
        CLKOUTB_EN      : string  := "TRUE";
        CLKOUTC_EN      : string  := "TRUE";
        CLKOUTD_EN      : string  := "TRUE";
        DYN_DTA_SEL     : string  := "FALSE";
        DYN_DTB_SEL     : string  := "FALSE";
        CLKOUTA_DT_DIR  : vl_logic := Hi1;
        CLKOUTB_DT_DIR  : vl_logic := Hi1;
        CLKOUTA_DT_STEP : integer := 0;
        CLKOUTB_DT_STEP : integer := 0;
        CLKA_IN_SEL     : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        CLKA_OUT_SEL    : vl_logic := Hi0;
        CLKB_IN_SEL     : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        CLKB_OUT_SEL    : vl_logic := Hi0;
        CLKC_IN_SEL     : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        CLKC_OUT_SEL    : vl_logic := Hi0;
        CLKD_IN_SEL     : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        CLKD_OUT_SEL    : vl_logic := Hi0;
        CLKFB_SEL       : string  := "INTERNAL";
        DYN_DPA_EN      : string  := "FALSE";
        DYN_PSB_SEL     : string  := "FALSE";
        DYN_PSC_SEL     : string  := "FALSE";
        DYN_PSD_SEL     : string  := "FALSE";
        PSB_COARSE      : integer := 1;
        PSB_FINE        : integer := 0;
        PSC_COARSE      : integer := 1;
        PSC_FINE        : integer := 0;
        PSD_COARSE      : integer := 1;
        PSD_FINE        : integer := 0;
        DTMS_ENB        : string  := "FALSE";
        DTMS_ENC        : string  := "FALSE";
        DTMS_END        : string  := "FALSE";
        RESET_I_EN      : string  := "FALSE";
        RESET_S_EN      : string  := "FALSE";
        DYN_ICP_SEL     : string  := "FALSE";
        ICP_SEL         : vl_logic_vector(0 to 4) := (HiX, HiX, HiX, HiX, HiX);
        DYN_RES_SEL     : string  := "FALSE";
        LPR_REF         : vl_logic_vector(0 to 6) := (HiX, HiX, HiX, HiX, HiX, HiX, HiX)
    );
    port(
        CLKOUTA         : out    vl_logic;
        CLKOUTB         : out    vl_logic;
        CLKOUTC         : out    vl_logic;
        CLKOUTD         : out    vl_logic;
        LOCK            : out    vl_logic;
        CLKIN           : in     vl_logic;
        CLKFB           : in     vl_logic;
        ENCLKA          : in     vl_logic;
        ENCLKB          : in     vl_logic;
        ENCLKC          : in     vl_logic;
        ENCLKD          : in     vl_logic;
        FBDSEL          : in     vl_logic_vector(5 downto 0);
        IDSEL           : in     vl_logic_vector(5 downto 0);
        ODSELA          : in     vl_logic_vector(6 downto 0);
        ODSELB          : in     vl_logic_vector(6 downto 0);
        ODSELC          : in     vl_logic_vector(6 downto 0);
        ODSELD          : in     vl_logic_vector(6 downto 0);
        DTA             : in     vl_logic_vector(3 downto 0);
        DTB             : in     vl_logic_vector(3 downto 0);
        PSSEL           : in     vl_logic_vector(1 downto 0);
        PSDIR           : in     vl_logic;
        PSPULSE         : in     vl_logic;
        ICPSEL          : in     vl_logic_vector(4 downto 0);
        LPFRES          : in     vl_logic_vector(2 downto 0);
        RESET           : in     vl_logic;
        RESET_P         : in     vl_logic;
        RESET_I         : in     vl_logic;
        RESET_S         : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of FCLKIN : constant is 1;
    attribute mti_svvh_generic_type of DYN_IDIV_SEL : constant is 1;
    attribute mti_svvh_generic_type of IDIV_SEL : constant is 1;
    attribute mti_svvh_generic_type of DYN_FBDIV_SEL : constant is 1;
    attribute mti_svvh_generic_type of FBDIV_SEL : constant is 1;
    attribute mti_svvh_generic_type of DYN_ODIVA_SEL : constant is 1;
    attribute mti_svvh_generic_type of ODIVA_SEL : constant is 1;
    attribute mti_svvh_generic_type of DYN_ODIVB_SEL : constant is 1;
    attribute mti_svvh_generic_type of ODIVB_SEL : constant is 1;
    attribute mti_svvh_generic_type of DYN_ODIVC_SEL : constant is 1;
    attribute mti_svvh_generic_type of ODIVC_SEL : constant is 1;
    attribute mti_svvh_generic_type of DYN_ODIVD_SEL : constant is 1;
    attribute mti_svvh_generic_type of ODIVD_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKOUTA_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUTB_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUTC_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUTD_EN : constant is 1;
    attribute mti_svvh_generic_type of DYN_DTA_SEL : constant is 1;
    attribute mti_svvh_generic_type of DYN_DTB_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKOUTA_DT_DIR : constant is 1;
    attribute mti_svvh_generic_type of CLKOUTB_DT_DIR : constant is 1;
    attribute mti_svvh_generic_type of CLKOUTA_DT_STEP : constant is 1;
    attribute mti_svvh_generic_type of CLKOUTB_DT_STEP : constant is 1;
    attribute mti_svvh_generic_type of CLKA_IN_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKA_OUT_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKB_IN_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKB_OUT_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKC_IN_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKC_OUT_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKD_IN_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKD_OUT_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKFB_SEL : constant is 1;
    attribute mti_svvh_generic_type of DYN_DPA_EN : constant is 1;
    attribute mti_svvh_generic_type of DYN_PSB_SEL : constant is 1;
    attribute mti_svvh_generic_type of DYN_PSC_SEL : constant is 1;
    attribute mti_svvh_generic_type of DYN_PSD_SEL : constant is 1;
    attribute mti_svvh_generic_type of PSB_COARSE : constant is 1;
    attribute mti_svvh_generic_type of PSB_FINE : constant is 1;
    attribute mti_svvh_generic_type of PSC_COARSE : constant is 1;
    attribute mti_svvh_generic_type of PSC_FINE : constant is 1;
    attribute mti_svvh_generic_type of PSD_COARSE : constant is 1;
    attribute mti_svvh_generic_type of PSD_FINE : constant is 1;
    attribute mti_svvh_generic_type of DTMS_ENB : constant is 1;
    attribute mti_svvh_generic_type of DTMS_ENC : constant is 1;
    attribute mti_svvh_generic_type of DTMS_END : constant is 1;
    attribute mti_svvh_generic_type of RESET_I_EN : constant is 1;
    attribute mti_svvh_generic_type of RESET_S_EN : constant is 1;
    attribute mti_svvh_generic_type of DYN_ICP_SEL : constant is 1;
    attribute mti_svvh_generic_type of ICP_SEL : constant is 1;
    attribute mti_svvh_generic_type of DYN_RES_SEL : constant is 1;
    attribute mti_svvh_generic_type of LPR_REF : constant is 1;
end PLLO;
